module random_generator(
    input wire clk,
    input wire rst_n,
    input wire load_seed,       // ��ư ���� �� High
    input wire [15:0] seed_val, // Top���� ��� ���� ī���� ��
    
    output reg [3:0] d1, // õ�� �ڸ�
    output reg [3:0] d2, // ���� �ڸ�
    output reg [3:0] d3, // ���� �ڸ�
    output reg [3:0] d4  // ���� �ڸ�
);

    reg [15:0] lfsr_reg;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            lfsr_reg <= 16'h1234; // �ʱⰪ
        end else if (load_seed) begin
            // �õ尪�� 0�̸� 1�� ���� ��ȯ (Lock-up ����)
            lfsr_reg <= (seed_val == 0) ? 16'h1 : seed_val;
        end else begin
            // 16-bit Galois LFSR
            lfsr_reg[15] <= lfsr_reg[14];
            lfsr_reg[14] <= lfsr_reg[13] ^ lfsr_reg[15];
            lfsr_reg[13] <= lfsr_reg[12] ^ lfsr_reg[15];
            lfsr_reg[12] <= lfsr_reg[11];
            lfsr_reg[11] <= lfsr_reg[10] ^ lfsr_reg[15];
            lfsr_reg[10] <= lfsr_reg[9];
            lfsr_reg[9:0] <= {lfsr_reg[8:0], lfsr_reg[15]};
        end
    end

    // ��� �й� (Combinational Logic)
    always @(*) begin
        d1 = lfsr_reg[15:12] % 10;
        d2 = lfsr_reg[11:8]  % 10;
        d3 = lfsr_reg[7:4]   % 10;
        d4 = lfsr_reg[3:0]   % 10;
    end
endmodule