module servo_controller(
    input clk,
    input rst,
    input [3:0] state,
    
    output reg servo // Servo motor�� �����ϱ� ���� pwm ��ȣ ���
);

localparam UNLOCK = 4'b0111; // �ݰ� ��� ���� state

localparam PWM_PERIOD = 1000000; // PWM�� �ֱ� (20ms)�� ���� ��ü ī��Ʈ ��

localparam DUTY_0_DEG = 50000; // 1.0ms pulse �� (���)
localparam DUTY_180_DEG = 100000; // 2.0ms pulse �� (����)

reg [19:0] pwm_counter;
reg [19:0] duty_cycle;

always @(posedge clk or posedge rst) begin
    if(rst) begin
        pwm_counter <= 20'd0;
        duty_cycle <= DUTY_0_DEG;
    end
    else begin
        if (pwm_counter == PWM_PERIOD-1) begin // 999,999���� ī���� ����
            pwm_counter <= 20'd0;
            
            // ���� state�� ���
            if(state == UNLOCK) begin
                duty_cycle <= DUTY_180_DEG; // ����
            end 
            // �� ���� state�� ���
            else begin
                duty_cycle <= DUTY_0_DEG; // ���
            end
        
        end else begin
            pwm_counter <= pwm_counter + 1;
        end
        
        // PWM Generation
        // �޽� �� �̳��� �� high ���
        if(pwm_counter < duty_cycle) begin
            servo <= 1'b1;
        end
        // �޽� �� �ʰ��ϸ� low ���
        else begin 
            servo <= 1'b0;
        end
    end
end

endmodule