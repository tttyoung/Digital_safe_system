module cal_result(
    // 1. ���� �Է� (4�ڸ�)
    input wire [3:0] d1, // õ�� �ڸ� (���� ����)
    input wire [3:0] d2,
    input wire [3:0] d3,
    input wire [3:0] d4, // ���� �ڸ� (���� ������)

    // 2. ������ �Է� (������ ��忡�� �� ��ȣ -> ������ ���Ƿ� ���� ����)
    input wire op1, // ù ��° ������ (d1 ? d2) : 0�̸� +, 1�̸� *
    input wire op2, // �� ��° ������ (Res ? d3)
    input wire op3, // �� ��° ������ (Res ? d4)

    // 3. ���� ���� ���
    output reg [15:0] correct_ans // �ִ� 9*9*9*9=6561 �̹Ƿ� 16��Ʈ�� ���
);

    // �߰� ��� ������ ������ ������
    // ������ ���̸� ���ڰ� Ŀ���Ƿ� �˳��ϰ� 16��Ʈ�� ����ϴ�.
    reg [15:0] step1_res; // (d1 op1 d2) ���
    reg [15:0] step2_res; // (step1 op2 d3) ���

    always @(*) begin
        // --- 1�ܰ�: d1�� d2 ���� ---
        if (op1 == 1'b0) step1_res = d1 + d2;      // ����
        else             step1_res = d1 * d2;      // ����

        // --- 2�ܰ�: 1�ܰ� ����� d3 ���� ---
        if (op2 == 1'b0) step2_res = step1_res + d3;
        else             step2_res = step1_res * d3;

        // --- 3�ܰ�: 2�ܰ� ����� d4 ���� (����) ---
        if (op3 == 1'b0) correct_ans = step2_res + d4;
        else             correct_ans = step2_res * d4;
    end

endmodule