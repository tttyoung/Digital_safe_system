module clock_divider(
    input clk,          // ���� �⺻ Ŭ�� (���� 50MHz)
    input rst_n,
    output reg clk_1khz, // 7-���׸�Ʈ ��ĵ�� (������ ������)
    output reg clk_1hz   // Ÿ�̸� ī��Ʈ�� (1��)
);
    // 50MHz = 50,000,000Hz
    // 1kHz�� ������� 50,000���� -> 25,000���� ���
    // 1Hz�� ������� 50,000,000���� -> 25,000,000���� ���
    
    integer cnt_1k = 0;
    integer cnt_1h = 0;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            cnt_1k <= 0; clk_1khz <= 0;
            cnt_1h <= 0; clk_1hz <= 0;
        end else begin
            // 1kHz ����
            if(cnt_1k >= 24999) begin // 50,000 / 2 - 1
                cnt_1k <= 0;
                clk_1khz <= ~clk_1khz;
            end else cnt_1k <= cnt_1k + 1;

            // 1Hz ����
            if(cnt_1h >= 24999999) begin // 50,000,000 / 2 - 1
                cnt_1h <= 0;
                clk_1hz <= ~clk_1hz;
            end else cnt_1h <= cnt_1h + 1;
        end
    end
endmodule