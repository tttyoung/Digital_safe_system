module adc_controller(
    input wire clk_500khz,   
    input wire rst_n,
    
    output wire adc_clk,     
    output reg adc_start,  // adc��ȯ���ۿ���  
    output reg adc_ale,    // adc_addr�� �Ƿ��ִ� ä�ι�ȣ ��ġ���ִ� ��ȣ
    output reg adc_oe,     // ��ȯ ����� ���������� 
    output reg [2:0] adc_addr, // adcä��
    input wire adc_eoc,  //��ȯ �� �Ǿ�����    
    input wire [7:0] adc_data_in,  //��ȯ��� 8��Ʈ ������
        
    // FSM �����
    output reg [7:0] dial_value // ���� ���(dial�� ���� ��)
);

    assign adc_clk = clk_500khz;

    // 2. �� ��Ű�� ���� (State Machine)
    reg [2:0] state;
    reg [7:0] wait_cnt; 

    localparam S_IDLE  = 0; // �غ�ܰ�
    localparam S_START = 1; // ��ɽ���
    localparam S_WAIT  = 2; // wait
    localparam S_READ  = 3; // ��� �б�

    // FSM�� 500kHz ���ڿ� ���缭 ����
    always @(posedge clk_500khz or negedge rst_n) begin
        if(!rst_n) begin
            state <= S_IDLE;
            adc_start <= 0; adc_ale <= 0; adc_oe <= 0;
            adc_addr <= 0; dial_value <= 0;
            wait_cnt <= 0;
        end else begin
            case(state)
                S_IDLE: begin //��� ��ȣ �ʱ�ȭ
                    adc_start <= 0; adc_ale <= 0; adc_oe <= 0;
                    state <= S_START;
                end
                
                S_START: begin
                    adc_addr <= 3'b000; // 0�� ä�� (��������)
                    adc_ale <= 1;       // �ּ� ��ġ
                    adc_start <= 1;     // ���� ��ȣ
                    state <= S_WAIT;
                    wait_cnt <= 0;
                end
                
                S_WAIT: begin
                    adc_ale <= 0;
                    adc_start <= 0;
                    
                    if(adc_eoc == 1 || wait_cnt > 60) begin 
                        state <= S_READ;
                    end else begin
                        wait_cnt <= wait_cnt + 1;
                    end
                end
                
                S_READ: begin
                    adc_oe <= 1; // ��� Ȱ��ȭ
                    dial_value <= adc_data_in; // ������ �б�
                    state <= S_IDLE;
                end
            endcase
        end
    end

endmodule