module timer(
    input wire clk,          
    input wire rst_n,        
    
    input wire clk_1hz,  //Ÿ�̸ӿ� 1hz Ŭ��    
    input wire run_timer,    //1: �ð����� ����
    input wire reset_timer,  //1: Ÿ�̸� �ٽ� 1������ ���½�Ű��
    
    // 0�̸� 1�� ���, 1�̸� 5�� ���
    input wire timer_mode_5min, 
    
    output reg [5:0] curr_min, 
    output reg [5:0] curr_sec, 
    output reg time_out    //�ð� ����    
);

    reg clk_1hz_prev;
    wire tick_1s;
    assign tick_1s = (clk_1hz == 1'b1) && (clk_1hz_prev == 1'b0);

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) clk_1hz_prev <= 0;
        else       clk_1hz_prev <= clk_1hz;
    end

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            curr_min <= 1; curr_sec <= 0; // �⺻ 1��
            time_out <= 0;
        end 
        else begin
            if (reset_timer) begin
                time_out <= 0;
                curr_sec <= 0;
                
                if (timer_mode_5min == 1'b1) 
                    curr_min <= 5; // ���� ���� 5��
                else 
                    curr_min <= 1; // ��ҿ��� 1��
            end 
            
            else if (run_timer && !time_out && tick_1s) begin
                if (curr_sec == 0) begin
                    if (curr_min == 0) begin
                        time_out <= 1; 
                    end else begin
                        curr_min <= curr_min - 1;
                        curr_sec <= 59;
                    end
                end else begin
                    curr_sec <= curr_sec - 1;
                end
            end
        end
    end

endmodule