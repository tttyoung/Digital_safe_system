module output_system_core(
    // �Է� ( FSM/��Ʈ�� �������� ���� ����)
    input clk, 
    input rst,
    input [3:0] state, // ���� FSM ����
    input [3:0] chance_count, // ���� ��ȸ ī��Ʈ
    input [15:0] input_data, // 8-7���׸�Ʈ�� ���� ��ǲ
    input [5:0] timer_min, // ����� minutes
    input [5:0] timer_sec, // ����� sec
    input clk_1khz, // PWM/Timing�� ���� 1KHZ clock
    input clk_mux, // 8-7���׸�Ʈ�� ���� ~500Hz Clock 
    
    // ���
    output [11:0] rgb_out, // FULL COLOR LED
    output [2:0] chance_led, // ���� ��ȸ led
    output servo_pwm, // servo motor
    output piezo, // piezo
    output[6:0] set_cathode, // 7���׸�Ʈ ���� ����� ����
    output[7:0] seg_anode, // 8-7���׸�Ʈ � �ڸ� ������� ����
    output[7:0] lcd_data, // text lcd
    output lcd_en, lcd_rs, lcd_rw // lcd ��Ʈ�ѿ� �ʿ��� ��ȣ
);

// wire ���� (��� ���� ��ȣ�� �����ϰų� �����͸� �ӽ÷� �����ϴµ� ���)
wire servo_pwm_out; // Servo Motor Controller ����� PWM ��� ��ȣ�� �ӽ÷� ����
wire [6:0] timer_seg_cathode_w; // ��⿡�� ������ 7���׸�Ʈ ���� �����͸� �ӽ÷� ���޹���
wire [7:0] timer_seg_anode_w; // ��⿡�� ������ 7���׸�Ʈ 8���� �� �ڸ� ��ȣ�� �ӽ÷� ����.

// ��� ��ü ����
// 1. feedback(FULL COLOR LED & Piezo)
feedback_controller U_FEEDBACK(
    .clk_1khz(clk_1khz),
    .rst(rst),
    .state(state),
    .rgb_out(rgb_out),
    .piezo_pwm(piezo_pwm)
);

// 2. �������� ��Ʈ�ѷ�

// 3. 8cell 7���׸�Ʈ display & chance led
timer_display_mux U_TIMER_DISPLAY(
    .clk_mux(clk_mux),
    .rst(rst),
    .state(state),
    .chance_count(chance_count),
    .input_data(input_data),
    .timer_min(timer_min),
    .timer_sec(timer_sec),
    .seg_cathode(seg_cathode), 
    .seg_anode(seg_anode),  
    .chance_led(chance_led)
);

// 4. �ؽ�Ʈ LCD
lcd_driver U_LCD (
    .clk(clk),
    .rst(rst),
    .state(state),
    .lcd_data(lcd_data),
    .lcd_en(lcd_en),
    .lcd_rs(lcd_rs),
    .lcd_rw(lcd_rw)
);

endmodule
