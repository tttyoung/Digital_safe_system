module keypad(
    input wire clk,          
    input wire rst_n,        
    
    // 0~9�� ��: ���� 0~9
    // 10�� ��: * (��)
    // 11�� ��: # (��)
    input wire [11:0] btn_in, //�������ڸ� 0   ex) 0���� ������ -> 111111111110
    
    output reg [3:0] key_value, // ���� ���� (0~15)
    output reg key_valid        // ���� ��ȣ (1 pulse)
);

    // ��ư ���� ������ ���� ��������
    reg [11:0] btn_prev;
    
    // 12�� ��ư �� �ϳ��� ���ȴ��� Ȯ��
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            btn_prev <= 12'hFFF; // ��� �� ���� ����(1)�� �ʱ�ȭ (�ʱⰪ: 111111111111)
            key_valid <= 0;
            key_value <= 0;
        end else begin
            btn_prev <= btn_in; // ���� ���� ������Ʈ(���� Ŭ�� ������)
            if (btn_prev != btn_in) begin              
                key_valid <= 1; // ������ȣ ����
                // � ��ư���� ã�� (�켱����: 0������ Ȯ��)
                if      (btn_prev[0] && !btn_in[0])  key_value <= 4'd0; // 0�� ��ư
                else if (btn_prev[1] && !btn_in[1])  key_value <= 4'd1; // 1�� ��ư
                else if (btn_prev[2] && !btn_in[2])  key_value <= 4'd2; // 2�� ��ư
                else if (btn_prev[3] && !btn_in[3])  key_value <= 4'd3; // 3�� ��ư
                else if (btn_prev[4] && !btn_in[4])  key_value <= 4'd4; // 4�� ��ư
                else if (btn_prev[5] && !btn_in[5])  key_value <= 4'd5; // 5�� ��ư
                else if (btn_prev[6] && !btn_in[6])  key_value <= 4'd6; // 6�� ��ư
                else if (btn_prev[7] && !btn_in[7])  key_value <= 4'd7; // 7�� ��ư
                else if (btn_prev[8] && !btn_in[8])  key_value <= 4'd8; // 8�� ��ư
                else if (btn_prev[9] && !btn_in[9])  key_value <= 4'd9; // 9�� ��ư
                else if (btn_prev[10] && !btn_in[10]) key_value <= 4'd14; // * (10�� ��)
                else if (btn_prev[11] && !btn_in[11]) key_value <= 4'd15; // # (11�� ��)
                else begin
                    // ���� �� �ƴ϶� ���� ���(0->1) ���� ����
                    key_valid <= 0; 
                end

            end else begin
                key_valid <= 0; // �ƹ� ��ȭ ����
            end
        end
    end

endmodule